module shiftRows_tb;

reg [127:0] in;
wire [127:0] out;	


shiftRows m (in,out);


initial begin
	$monitor("input= %H , output= %h",in,out);
	in = 128'hd42711aee0bf98f1b8b45de51e415230;
end
endmodule